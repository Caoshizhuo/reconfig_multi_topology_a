library verilog;
use verilog.vl_types.all;
entity reconfig_multi_topology_a_tb is
end reconfig_multi_topology_a_tb;
